`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:00:24 07/05/2016 
// Design Name: 
// Module Name:    exp_adjust
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module add(
    input [4:0] a,
    input [4:0] exp_adjust,
    output [5:0] c
    );

assign c = a - exp_adjust ;

endmodule
